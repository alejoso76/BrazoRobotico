`timescale 1ns / 1ps
//-------------------------------------------------------------------

module memoriaRAM(
    input CLK,
    input [7:0] address,
	 input [31:0] data,
    output reg [31:0] DATOS
    );

//-------------------------------------------------------------------
always @(posedge CLK)
	begin                   
		
	end
endmodule
